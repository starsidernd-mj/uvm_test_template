`ifndef COVERAGE_SVH
`define COVERAGE_SVH

import uvm_pkg::*;

`include "uvm_macros.svh"

`endif
