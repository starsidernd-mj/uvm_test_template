`ifndef GEN_ITEM_SEQ_SVH
`define GEN_ITEM_SEQ_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`include "Item.sv"

`endif
