`ifndef MONITOR_SVH
`define MONITOR_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`include "../../env/sequencers/Item.sv"

`endif
