`ifndef BASE_TEST_SVH
`define BASE_TEST_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../my_macros.svh"

`include "../env/env.sv"
`include "../env/sequencers/gen_item_seq.sv"

`endif
