`ifndef SCOREBOARD_SVH
`define SCOREBOARD_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`include "../sequencers/Item.sv"

`endif
