`ifndef MY_MACROS_SVH
`define MY_MACROS_SVH

`define LENGTH 4



`endif
