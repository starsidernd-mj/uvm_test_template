`ifndef DES_IF_SVH
`define DES_IF_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`endif
