`ifndef ITEM_SVH
`define ITEM_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`endif
