`ifndef TEST_1011_SVH
`define TEST_1011_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../my_macros.svh"
`include "../env/env.sv"
`include "base_test.sv"
`include "../env/sequencers/gen_item_seq.sv"

`endif
