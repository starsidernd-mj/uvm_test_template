`ifndef DRIVER_SVH
`define DRIVER_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`include "../../env/sequencers/Item.sv"

`endif
