`ifndef COVERAGE_VIF_SVH
`define COVERAGE_VIF_SVH

//include the UVM package
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "../../my_macros.svh"

`endif

